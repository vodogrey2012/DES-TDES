`timescale 1ns/10ps

module f
    (
    input [31:0] R,
    input [31:0] L,
    input [47:0] k,
    output logic [31:0] R_out,
    output logic [31:0] L_out
    );

assign L_out = R;

// E permutation
logic [47:0] R_ext;
assign R_ext = {R[0],  R[31], R[30], R[29], R[28], R[27], 
                R[28], R[27], R[26], R[25], R[24], R[23],
                R[24], R[23], R[22], R[21], R[20], R[19],
                R[20], R[19], R[18], R[17], R[16], R[15],
                R[16], R[15], R[14], R[13], R[12], R[11],
                R[12], R[11], R[10], R[9],  R[8],  R[7],
                R[8],  R[7],  R[6],  R[5],  R[4],  R[3],
                R[4],  R[3],  R[2],  R[1],  R[0],  R[31]};

// xor with key
logic [47:0] xor_result;
assign xor_result = R_ext ^ k;

// S calculation
logic [31:0] S;

always_comb
begin
    case ({xor_result[47], xor_result[42], xor_result[46:43]})
        {2'd0, 4'd0}:  S[31:28] = 4'd14;
        {2'd0, 4'd1}:  S[31:28] = 4'd4;
        {2'd0, 4'd2}:  S[31:28] = 4'd13;
        {2'd0, 4'd3}:  S[31:28] = 4'd1;
        {2'd0, 4'd4}:  S[31:28] = 4'd2;
        {2'd0, 4'd5}:  S[31:28] = 4'd15;
        {2'd0, 4'd6}:  S[31:28] = 4'd11;
        {2'd0, 4'd7}:  S[31:28] = 4'd8;
        {2'd0, 4'd8}:  S[31:28] = 4'd3;
        {2'd0, 4'd9}:  S[31:28] = 4'd10;
        {2'd0, 4'd10}: S[31:28] = 4'd6;
        {2'd0, 4'd11}: S[31:28] = 4'd12;
        {2'd0, 4'd12}: S[31:28] = 4'd5;
        {2'd0, 4'd13}: S[31:28] = 4'd9;
        {2'd0, 4'd14}: S[31:28] = 4'd0;
        {2'd0, 4'd15}: S[31:28] = 4'd7;
        {2'd1, 4'd0}:  S[31:28] = 4'd0;
        {2'd1, 4'd1}:  S[31:28] = 4'd15;
        {2'd1, 4'd2}:  S[31:28] = 4'd7;
        {2'd1, 4'd3}:  S[31:28] = 4'd4;
        {2'd1, 4'd4}:  S[31:28] = 4'd14;
        {2'd1, 4'd5}:  S[31:28] = 4'd2;
        {2'd1, 4'd6}:  S[31:28] = 4'd13;
        {2'd1, 4'd7}:  S[31:28] = 4'd1;
        {2'd1, 4'd8}:  S[31:28] = 4'd10;
        {2'd1, 4'd9}:  S[31:28] = 4'd6;
        {2'd1, 4'd10}: S[31:28] = 4'd12;
        {2'd1, 4'd11}: S[31:28] = 4'd11;
        {2'd1, 4'd12}: S[31:28] = 4'd9;
        {2'd1, 4'd13}: S[31:28] = 4'd5;
        {2'd1, 4'd14}: S[31:28] = 4'd3;
        {2'd1, 4'd15}: S[31:28] = 4'd8;
        {2'd2, 4'd0}:  S[31:28] = 4'd4;
        {2'd2, 4'd1}:  S[31:28] = 4'd1;
        {2'd2, 4'd2}:  S[31:28] = 4'd14;
        {2'd2, 4'd3}:  S[31:28] = 4'd8;
        {2'd2, 4'd4}:  S[31:28] = 4'd13;
        {2'd2, 4'd5}:  S[31:28] = 4'd6;
        {2'd2, 4'd6}:  S[31:28] = 4'd2;
        {2'd2, 4'd7}:  S[31:28] = 4'd11;
        {2'd2, 4'd8}:  S[31:28] = 4'd15;
        {2'd2, 4'd9}:  S[31:28] = 4'd12;
        {2'd2, 4'd10}: S[31:28] = 4'd9;
        {2'd2, 4'd11}: S[31:28] = 4'd7;
        {2'd2, 4'd12}: S[31:28] = 4'd3;
        {2'd2, 4'd13}: S[31:28] = 4'd10;
        {2'd2, 4'd14}: S[31:28] = 4'd5;
        {2'd2, 4'd15}: S[31:28] = 4'd0;
        {2'd3, 4'd0}:  S[31:28] = 4'd15;
        {2'd3, 4'd1}:  S[31:28] = 4'd12;
        {2'd3, 4'd2}:  S[31:28] = 4'd8;
        {2'd3, 4'd3}:  S[31:28] = 4'd2;
        {2'd3, 4'd4}:  S[31:28] = 4'd4;
        {2'd3, 4'd5}:  S[31:28] = 4'd9;
        {2'd3, 4'd6}:  S[31:28] = 4'd1;
        {2'd3, 4'd7}:  S[31:28] = 4'd7;
        {2'd3, 4'd8}:  S[31:28] = 4'd5;
        {2'd3, 4'd9}:  S[31:28] = 4'd11;
        {2'd3, 4'd10}: S[31:28] = 4'd3;
        {2'd3, 4'd11}: S[31:28] = 4'd14;
        {2'd3, 4'd12}: S[31:28] = 4'd10;
        {2'd3, 4'd13}: S[31:28] = 4'd0;
        {2'd3, 4'd14}: S[31:28] = 4'd6;
        {2'd3, 4'd15}: S[31:28] = 4'd13;
endcase
end

always_comb
begin
    case ({xor_result[41], xor_result[36], xor_result[40:37]})
        {2'd0, 4'd0}:  S[27:24] = 4'd15;
        {2'd0, 4'd1}:  S[27:24] = 4'd1;
        {2'd0, 4'd2}:  S[27:24] = 4'd8;
        {2'd0, 4'd3}:  S[27:24] = 4'd14;
        {2'd0, 4'd4}:  S[27:24] = 4'd6;
        {2'd0, 4'd5}:  S[27:24] = 4'd11;
        {2'd0, 4'd6}:  S[27:24] = 4'd3;
        {2'd0, 4'd7}:  S[27:24] = 4'd4;
        {2'd0, 4'd8}:  S[27:24] = 4'd9;
        {2'd0, 4'd9}:  S[27:24] = 4'd7;
        {2'd0, 4'd10}: S[27:24] = 4'd2;
        {2'd0, 4'd11}: S[27:24] = 4'd13;
        {2'd0, 4'd12}: S[27:24] = 4'd12;
        {2'd0, 4'd13}: S[27:24] = 4'd0;
        {2'd0, 4'd14}: S[27:24] = 4'd5;
        {2'd0, 4'd15}: S[27:24] = 4'd10;
        {2'd1, 4'd0}:  S[27:24] = 4'd3;
        {2'd1, 4'd1}:  S[27:24] = 4'd13;
        {2'd1, 4'd2}:  S[27:24] = 4'd4;
        {2'd1, 4'd3}:  S[27:24] = 4'd7;
        {2'd1, 4'd4}:  S[27:24] = 4'd15;
        {2'd1, 4'd5}:  S[27:24] = 4'd2;
        {2'd1, 4'd6}:  S[27:24] = 4'd8;
        {2'd1, 4'd7}:  S[27:24] = 4'd14;
        {2'd1, 4'd8}:  S[27:24] = 4'd12;
        {2'd1, 4'd9}:  S[27:24] = 4'd0;
        {2'd1, 4'd10}: S[27:24] = 4'd1;
        {2'd1, 4'd11}: S[27:24] = 4'd10;
        {2'd1, 4'd12}: S[27:24] = 4'd6;
        {2'd1, 4'd13}: S[27:24] = 4'd9;
        {2'd1, 4'd14}: S[27:24] = 4'd11;
        {2'd1, 4'd15}: S[27:24] = 4'd5;
        {2'd2, 4'd0}:  S[27:24] = 4'd0;
        {2'd2, 4'd1}:  S[27:24] = 4'd14;
        {2'd2, 4'd2}:  S[27:24] = 4'd7;
        {2'd2, 4'd3}:  S[27:24] = 4'd11;
        {2'd2, 4'd4}:  S[27:24] = 4'd10;
        {2'd2, 4'd5}:  S[27:24] = 4'd4;
        {2'd2, 4'd6}:  S[27:24] = 4'd13;
        {2'd2, 4'd7}:  S[27:24] = 4'd1;
        {2'd2, 4'd8}:  S[27:24] = 4'd5;
        {2'd2, 4'd9}:  S[27:24] = 4'd8;
        {2'd2, 4'd10}: S[27:24] = 4'd12;
        {2'd2, 4'd11}: S[27:24] = 4'd6;
        {2'd2, 4'd12}: S[27:24] = 4'd9;
        {2'd2, 4'd13}: S[27:24] = 4'd3;
        {2'd2, 4'd14}: S[27:24] = 4'd2;
        {2'd2, 4'd15}: S[27:24] = 4'd15;
        {2'd3, 4'd0}:  S[27:24] = 4'd13;
        {2'd3, 4'd1}:  S[27:24] = 4'd8;
        {2'd3, 4'd2}:  S[27:24] = 4'd10;
        {2'd3, 4'd3}:  S[27:24] = 4'd1;
        {2'd3, 4'd4}:  S[27:24] = 4'd3;
        {2'd3, 4'd5}:  S[27:24] = 4'd15;
        {2'd3, 4'd6}:  S[27:24] = 4'd4;
        {2'd3, 4'd7}:  S[27:24] = 4'd2;
        {2'd3, 4'd8}:  S[27:24] = 4'd11;
        {2'd3, 4'd9}:  S[27:24] = 4'd6;
        {2'd3, 4'd10}: S[27:24] = 4'd7;
        {2'd3, 4'd11}: S[27:24] = 4'd12;
        {2'd3, 4'd12}: S[27:24] = 4'd0;
        {2'd3, 4'd13}: S[27:24] = 4'd5;
        {2'd3, 4'd14}: S[27:24] = 4'd14;
        {2'd3, 4'd15}: S[27:24] = 4'd9;
endcase
end

always_comb
begin
    case ({xor_result[35], xor_result[30], xor_result[34:31]})
        {2'd0, 4'd0}:  S[23:20] = 4'd10;
        {2'd0, 4'd1}:  S[23:20] = 4'd0;
        {2'd0, 4'd2}:  S[23:20] = 4'd9;
        {2'd0, 4'd3}:  S[23:20] = 4'd14;
        {2'd0, 4'd4}:  S[23:20] = 4'd6;
        {2'd0, 4'd5}:  S[23:20] = 4'd3;
        {2'd0, 4'd6}:  S[23:20] = 4'd15;
        {2'd0, 4'd7}:  S[23:20] = 4'd5;
        {2'd0, 4'd8}:  S[23:20] = 4'd1;
        {2'd0, 4'd9}:  S[23:20] = 4'd13;
        {2'd0, 4'd10}: S[23:20] = 4'd12;
        {2'd0, 4'd11}: S[23:20] = 4'd7;
        {2'd0, 4'd12}: S[23:20] = 4'd11;
        {2'd0, 4'd13}: S[23:20] = 4'd4;
        {2'd0, 4'd14}: S[23:20] = 4'd2;
        {2'd0, 4'd15}: S[23:20] = 4'd8;
        {2'd1, 4'd0}:  S[23:20] = 4'd13;
        {2'd1, 4'd1}:  S[23:20] = 4'd7;
        {2'd1, 4'd2}:  S[23:20] = 4'd0;
        {2'd1, 4'd3}:  S[23:20] = 4'd9;
        {2'd1, 4'd4}:  S[23:20] = 4'd3;
        {2'd1, 4'd5}:  S[23:20] = 4'd4;
        {2'd1, 4'd6}:  S[23:20] = 4'd6;
        {2'd1, 4'd7}:  S[23:20] = 4'd10;
        {2'd1, 4'd8}:  S[23:20] = 4'd2;
        {2'd1, 4'd9}:  S[23:20] = 4'd8;
        {2'd1, 4'd10}: S[23:20] = 4'd5;
        {2'd1, 4'd11}: S[23:20] = 4'd14;
        {2'd1, 4'd12}: S[23:20] = 4'd12;
        {2'd1, 4'd13}: S[23:20] = 4'd11;
        {2'd1, 4'd14}: S[23:20] = 4'd15;
        {2'd1, 4'd15}: S[23:20] = 4'd1;
        {2'd2, 4'd0}:  S[23:20] = 4'd13;
        {2'd2, 4'd1}:  S[23:20] = 4'd6;
        {2'd2, 4'd2}:  S[23:20] = 4'd4;
        {2'd2, 4'd3}:  S[23:20] = 4'd9;
        {2'd2, 4'd4}:  S[23:20] = 4'd8;
        {2'd2, 4'd5}:  S[23:20] = 4'd15;
        {2'd2, 4'd6}:  S[23:20] = 4'd3;
        {2'd2, 4'd7}:  S[23:20] = 4'd0;
        {2'd2, 4'd8}:  S[23:20] = 4'd11;
        {2'd2, 4'd9}:  S[23:20] = 4'd1;
        {2'd2, 4'd10}: S[23:20] = 4'd2;
        {2'd2, 4'd11}: S[23:20] = 4'd12;
        {2'd2, 4'd12}: S[23:20] = 4'd5;
        {2'd2, 4'd13}: S[23:20] = 4'd10;
        {2'd2, 4'd14}: S[23:20] = 4'd14;
        {2'd2, 4'd15}: S[23:20] = 4'd7;
        {2'd3, 4'd0}:  S[23:20] = 4'd1;
        {2'd3, 4'd1}:  S[23:20] = 4'd10;
        {2'd3, 4'd2}:  S[23:20] = 4'd13;
        {2'd3, 4'd3}:  S[23:20] = 4'd0;
        {2'd3, 4'd4}:  S[23:20] = 4'd6;
        {2'd3, 4'd5}:  S[23:20] = 4'd9;
        {2'd3, 4'd6}:  S[23:20] = 4'd8;
        {2'd3, 4'd7}:  S[23:20] = 4'd7;
        {2'd3, 4'd8}:  S[23:20] = 4'd4;
        {2'd3, 4'd9}:  S[23:20] = 4'd15;
        {2'd3, 4'd10}: S[23:20] = 4'd14;
        {2'd3, 4'd11}: S[23:20] = 4'd3;
        {2'd3, 4'd12}: S[23:20] = 4'd11;
        {2'd3, 4'd13}: S[23:20] = 4'd5;
        {2'd3, 4'd14}: S[23:20] = 4'd2;
        {2'd3, 4'd15}: S[23:20] = 4'd12;
endcase
end

always_comb
begin
    case ({xor_result[29], xor_result[24], xor_result[28:25]})
        {2'd0, 4'd0}:  S[19:16] = 4'd7;
        {2'd0, 4'd1}:  S[19:16] = 4'd13;
        {2'd0, 4'd2}:  S[19:16] = 4'd14;
        {2'd0, 4'd3}:  S[19:16] = 4'd3;
        {2'd0, 4'd4}:  S[19:16] = 4'd0;
        {2'd0, 4'd5}:  S[19:16] = 4'd6;
        {2'd0, 4'd6}:  S[19:16] = 4'd9;
        {2'd0, 4'd7}:  S[19:16] = 4'd10;
        {2'd0, 4'd8}:  S[19:16] = 4'd1;
        {2'd0, 4'd9}:  S[19:16] = 4'd2;
        {2'd0, 4'd10}: S[19:16] = 4'd8;
        {2'd0, 4'd11}: S[19:16] = 4'd5;
        {2'd0, 4'd12}: S[19:16] = 4'd11;
        {2'd0, 4'd13}: S[19:16] = 4'd12;
        {2'd0, 4'd14}: S[19:16] = 4'd4;
        {2'd0, 4'd15}: S[19:16] = 4'd15;
        {2'd1, 4'd0}:  S[19:16] = 4'd13;
        {2'd1, 4'd1}:  S[19:16] = 4'd8;
        {2'd1, 4'd2}:  S[19:16] = 4'd11;
        {2'd1, 4'd3}:  S[19:16] = 4'd5;
        {2'd1, 4'd4}:  S[19:16] = 4'd6;
        {2'd1, 4'd5}:  S[19:16] = 4'd15;
        {2'd1, 4'd6}:  S[19:16] = 4'd0;
        {2'd1, 4'd7}:  S[19:16] = 4'd3;
        {2'd1, 4'd8}:  S[19:16] = 4'd4;
        {2'd1, 4'd9}:  S[19:16] = 4'd7;
        {2'd1, 4'd10}: S[19:16] = 4'd2;
        {2'd1, 4'd11}: S[19:16] = 4'd12;
        {2'd1, 4'd12}: S[19:16] = 4'd1;
        {2'd1, 4'd13}: S[19:16] = 4'd10;
        {2'd1, 4'd14}: S[19:16] = 4'd14;
        {2'd1, 4'd15}: S[19:16] = 4'd9;
        {2'd2, 4'd0}:  S[19:16] = 4'd10;
        {2'd2, 4'd1}:  S[19:16] = 4'd6;
        {2'd2, 4'd2}:  S[19:16] = 4'd9;
        {2'd2, 4'd3}:  S[19:16] = 4'd0;
        {2'd2, 4'd4}:  S[19:16] = 4'd12;
        {2'd2, 4'd5}:  S[19:16] = 4'd11;
        {2'd2, 4'd6}:  S[19:16] = 4'd7;
        {2'd2, 4'd7}:  S[19:16] = 4'd13;
        {2'd2, 4'd8}:  S[19:16] = 4'd15;
        {2'd2, 4'd9}:  S[19:16] = 4'd1;
        {2'd2, 4'd10}: S[19:16] = 4'd3;
        {2'd2, 4'd11}: S[19:16] = 4'd14;
        {2'd2, 4'd12}: S[19:16] = 4'd5;
        {2'd2, 4'd13}: S[19:16] = 4'd2;
        {2'd2, 4'd14}: S[19:16] = 4'd8;
        {2'd2, 4'd15}: S[19:16] = 4'd4;
        {2'd3, 4'd0}:  S[19:16] = 4'd3;
        {2'd3, 4'd1}:  S[19:16] = 4'd15;
        {2'd3, 4'd2}:  S[19:16] = 4'd0;
        {2'd3, 4'd3}:  S[19:16] = 4'd6;
        {2'd3, 4'd4}:  S[19:16] = 4'd10;
        {2'd3, 4'd5}:  S[19:16] = 4'd1;
        {2'd3, 4'd6}:  S[19:16] = 4'd13;
        {2'd3, 4'd7}:  S[19:16] = 4'd8;
        {2'd3, 4'd8}:  S[19:16] = 4'd9;
        {2'd3, 4'd9}:  S[19:16] = 4'd4;
        {2'd3, 4'd10}: S[19:16] = 4'd5;
        {2'd3, 4'd11}: S[19:16] = 4'd11;
        {2'd3, 4'd12}: S[19:16] = 4'd12;
        {2'd3, 4'd13}: S[19:16] = 4'd7;
        {2'd3, 4'd14}: S[19:16] = 4'd2;
        {2'd3, 4'd15}: S[19:16] = 4'd14;
endcase
end

always_comb
begin
    case ({xor_result[23], xor_result[18], xor_result[22:19]})
        {2'd0, 4'd0}:  S[15:12] = 4'd2;
        {2'd0, 4'd1}:  S[15:12] = 4'd12;
        {2'd0, 4'd2}:  S[15:12] = 4'd4;
        {2'd0, 4'd3}:  S[15:12] = 4'd1;
        {2'd0, 4'd4}:  S[15:12] = 4'd7;
        {2'd0, 4'd5}:  S[15:12] = 4'd10;
        {2'd0, 4'd6}:  S[15:12] = 4'd11;
        {2'd0, 4'd7}:  S[15:12] = 4'd6;
        {2'd0, 4'd8}:  S[15:12] = 4'd8;
        {2'd0, 4'd9}:  S[15:12] = 4'd5;
        {2'd0, 4'd10}: S[15:12] = 4'd3;
        {2'd0, 4'd11}: S[15:12] = 4'd15;
        {2'd0, 4'd12}: S[15:12] = 4'd13;
        {2'd0, 4'd13}: S[15:12] = 4'd0;
        {2'd0, 4'd14}: S[15:12] = 4'd14;
        {2'd0, 4'd15}: S[15:12] = 4'd9;
        {2'd1, 4'd0}:  S[15:12] = 4'd14;
        {2'd1, 4'd1}:  S[15:12] = 4'd11;
        {2'd1, 4'd2}:  S[15:12] = 4'd2;
        {2'd1, 4'd3}:  S[15:12] = 4'd12;
        {2'd1, 4'd4}:  S[15:12] = 4'd4;
        {2'd1, 4'd5}:  S[15:12] = 4'd7;
        {2'd1, 4'd6}:  S[15:12] = 4'd13;
        {2'd1, 4'd7}:  S[15:12] = 4'd1;
        {2'd1, 4'd8}:  S[15:12] = 4'd5;
        {2'd1, 4'd9}:  S[15:12] = 4'd0;
        {2'd1, 4'd10}: S[15:12] = 4'd15;
        {2'd1, 4'd11}: S[15:12] = 4'd10;
        {2'd1, 4'd12}: S[15:12] = 4'd3;
        {2'd1, 4'd13}: S[15:12] = 4'd9;
        {2'd1, 4'd14}: S[15:12] = 4'd8;
        {2'd1, 4'd15}: S[15:12] = 4'd6;
        {2'd2, 4'd0}:  S[15:12] = 4'd4;
        {2'd2, 4'd1}:  S[15:12] = 4'd2;
        {2'd2, 4'd2}:  S[15:12] = 4'd1;
        {2'd2, 4'd3}:  S[15:12] = 4'd11;
        {2'd2, 4'd4}:  S[15:12] = 4'd10;
        {2'd2, 4'd5}:  S[15:12] = 4'd13;
        {2'd2, 4'd6}:  S[15:12] = 4'd7;
        {2'd2, 4'd7}:  S[15:12] = 4'd8;
        {2'd2, 4'd8}:  S[15:12] = 4'd15;
        {2'd2, 4'd9}:  S[15:12] = 4'd9;
        {2'd2, 4'd10}: S[15:12] = 4'd12;
        {2'd2, 4'd11}: S[15:12] = 4'd5;
        {2'd2, 4'd12}: S[15:12] = 4'd6;
        {2'd2, 4'd13}: S[15:12] = 4'd3;
        {2'd2, 4'd14}: S[15:12] = 4'd0;
        {2'd2, 4'd15}: S[15:12] = 4'd14;
        {2'd3, 4'd0}:  S[15:12] = 4'd11;
        {2'd3, 4'd1}:  S[15:12] = 4'd8;
        {2'd3, 4'd2}:  S[15:12] = 4'd12;
        {2'd3, 4'd3}:  S[15:12] = 4'd7;
        {2'd3, 4'd4}:  S[15:12] = 4'd1;
        {2'd3, 4'd5}:  S[15:12] = 4'd14;
        {2'd3, 4'd6}:  S[15:12] = 4'd2;
        {2'd3, 4'd7}:  S[15:12] = 4'd13;
        {2'd3, 4'd8}:  S[15:12] = 4'd6;
        {2'd3, 4'd9}:  S[15:12] = 4'd15;
        {2'd3, 4'd10}: S[15:12] = 4'd0;
        {2'd3, 4'd11}: S[15:12] = 4'd9;
        {2'd3, 4'd12}: S[15:12] = 4'd10;
        {2'd3, 4'd13}: S[15:12] = 4'd4;
        {2'd3, 4'd14}: S[15:12] = 4'd5;
        {2'd3, 4'd15}: S[15:12] = 4'd3;
endcase
end

always_comb
begin
    case ({xor_result[17], xor_result[12], xor_result[16:13]})
        {2'd0, 4'd0}:  S[11:8] = 4'd12;
        {2'd0, 4'd1}:  S[11:8] = 4'd1;
        {2'd0, 4'd2}:  S[11:8] = 4'd10;
        {2'd0, 4'd3}:  S[11:8] = 4'd15;
        {2'd0, 4'd4}:  S[11:8] = 4'd9;
        {2'd0, 4'd5}:  S[11:8] = 4'd2;
        {2'd0, 4'd6}:  S[11:8] = 4'd6;
        {2'd0, 4'd7}:  S[11:8] = 4'd8;
        {2'd0, 4'd8}:  S[11:8] = 4'd0;
        {2'd0, 4'd9}:  S[11:8] = 4'd13;
        {2'd0, 4'd10}: S[11:8] = 4'd3;
        {2'd0, 4'd11}: S[11:8] = 4'd4;
        {2'd0, 4'd12}: S[11:8] = 4'd14;
        {2'd0, 4'd13}: S[11:8] = 4'd7;
        {2'd0, 4'd14}: S[11:8] = 4'd5;
        {2'd0, 4'd15}: S[11:8] = 4'd11;
        {2'd1, 4'd0}:  S[11:8] = 4'd10;
        {2'd1, 4'd1}:  S[11:8] = 4'd15;
        {2'd1, 4'd2}:  S[11:8] = 4'd4;
        {2'd1, 4'd3}:  S[11:8] = 4'd2;
        {2'd1, 4'd4}:  S[11:8] = 4'd7;
        {2'd1, 4'd5}:  S[11:8] = 4'd12;
        {2'd1, 4'd6}:  S[11:8] = 4'd9;
        {2'd1, 4'd7}:  S[11:8] = 4'd5;
        {2'd1, 4'd8}:  S[11:8] = 4'd6;
        {2'd1, 4'd9}:  S[11:8] = 4'd1;
        {2'd1, 4'd10}: S[11:8] = 4'd13;
        {2'd1, 4'd11}: S[11:8] = 4'd14;
        {2'd1, 4'd12}: S[11:8] = 4'd0;
        {2'd1, 4'd13}: S[11:8] = 4'd11;
        {2'd1, 4'd14}: S[11:8] = 4'd3;
        {2'd1, 4'd15}: S[11:8] = 4'd8;
        {2'd2, 4'd0}:  S[11:8] = 4'd9;
        {2'd2, 4'd1}:  S[11:8] = 4'd14;
        {2'd2, 4'd2}:  S[11:8] = 4'd15;
        {2'd2, 4'd3}:  S[11:8] = 4'd5;
        {2'd2, 4'd4}:  S[11:8] = 4'd2;
        {2'd2, 4'd5}:  S[11:8] = 4'd8;
        {2'd2, 4'd6}:  S[11:8] = 4'd12;
        {2'd2, 4'd7}:  S[11:8] = 4'd3;
        {2'd2, 4'd8}:  S[11:8] = 4'd7;
        {2'd2, 4'd9}:  S[11:8] = 4'd0;
        {2'd2, 4'd10}: S[11:8] = 4'd4;
        {2'd2, 4'd11}: S[11:8] = 4'd10;
        {2'd2, 4'd12}: S[11:8] = 4'd1;
        {2'd2, 4'd13}: S[11:8] = 4'd13;
        {2'd2, 4'd14}: S[11:8] = 4'd11;
        {2'd2, 4'd15}: S[11:8] = 4'd6;
        {2'd3, 4'd0}:  S[11:8] = 4'd4;
        {2'd3, 4'd1}:  S[11:8] = 4'd3;
        {2'd3, 4'd2}:  S[11:8] = 4'd2;
        {2'd3, 4'd3}:  S[11:8] = 4'd12;
        {2'd3, 4'd4}:  S[11:8] = 4'd9;
        {2'd3, 4'd5}:  S[11:8] = 4'd5;
        {2'd3, 4'd6}:  S[11:8] = 4'd15;
        {2'd3, 4'd7}:  S[11:8] = 4'd10;
        {2'd3, 4'd8}:  S[11:8] = 4'd11;
        {2'd3, 4'd9}:  S[11:8] = 4'd14;
        {2'd3, 4'd10}: S[11:8] = 4'd1;
        {2'd3, 4'd11}: S[11:8] = 4'd7;
        {2'd3, 4'd12}: S[11:8] = 4'd6;
        {2'd3, 4'd13}: S[11:8] = 4'd0;
        {2'd3, 4'd14}: S[11:8] = 4'd8;
        {2'd3, 4'd15}: S[11:8] = 4'd13;
endcase
end

always_comb
begin
    case ({xor_result[11], xor_result[6], xor_result[10:7]})
        {2'd0, 4'd0}:  S[7:4] = 4'd4;
        {2'd0, 4'd1}:  S[7:4] = 4'd11;
        {2'd0, 4'd2}:  S[7:4] = 4'd2;
        {2'd0, 4'd3}:  S[7:4] = 4'd14;
        {2'd0, 4'd4}:  S[7:4] = 4'd15;
        {2'd0, 4'd5}:  S[7:4] = 4'd0;
        {2'd0, 4'd6}:  S[7:4] = 4'd8;
        {2'd0, 4'd7}:  S[7:4] = 4'd13;
        {2'd0, 4'd8}:  S[7:4] = 4'd3;
        {2'd0, 4'd9}:  S[7:4] = 4'd12;
        {2'd0, 4'd10}: S[7:4] = 4'd9;
        {2'd0, 4'd11}: S[7:4] = 4'd7;
        {2'd0, 4'd12}: S[7:4] = 4'd5;
        {2'd0, 4'd13}: S[7:4] = 4'd10;
        {2'd0, 4'd14}: S[7:4] = 4'd6;
        {2'd0, 4'd15}: S[7:4] = 4'd1;
        {2'd1, 4'd0}:  S[7:4] = 4'd13;
        {2'd1, 4'd1}:  S[7:4] = 4'd0;
        {2'd1, 4'd2}:  S[7:4] = 4'd11;
        {2'd1, 4'd3}:  S[7:4] = 4'd7;
        {2'd1, 4'd4}:  S[7:4] = 4'd4;
        {2'd1, 4'd5}:  S[7:4] = 4'd9;
        {2'd1, 4'd6}:  S[7:4] = 4'd1;
        {2'd1, 4'd7}:  S[7:4] = 4'd10;
        {2'd1, 4'd8}:  S[7:4] = 4'd14;
        {2'd1, 4'd9}:  S[7:4] = 4'd3;
        {2'd1, 4'd10}: S[7:4] = 4'd5;
        {2'd1, 4'd11}: S[7:4] = 4'd12;
        {2'd1, 4'd12}: S[7:4] = 4'd2;
        {2'd1, 4'd13}: S[7:4] = 4'd15;
        {2'd1, 4'd14}: S[7:4] = 4'd8;
        {2'd1, 4'd15}: S[7:4] = 4'd6;
        {2'd2, 4'd0}:  S[7:4] = 4'd1;
        {2'd2, 4'd1}:  S[7:4] = 4'd4;
        {2'd2, 4'd2}:  S[7:4] = 4'd11;
        {2'd2, 4'd3}:  S[7:4] = 4'd13;
        {2'd2, 4'd4}:  S[7:4] = 4'd12;
        {2'd2, 4'd5}:  S[7:4] = 4'd3;
        {2'd2, 4'd6}:  S[7:4] = 4'd7;
        {2'd2, 4'd7}:  S[7:4] = 4'd14;
        {2'd2, 4'd8}:  S[7:4] = 4'd10;
        {2'd2, 4'd9}:  S[7:4] = 4'd15;
        {2'd2, 4'd10}: S[7:4] = 4'd6;
        {2'd2, 4'd11}: S[7:4] = 4'd8;
        {2'd2, 4'd12}: S[7:4] = 4'd0;
        {2'd2, 4'd13}: S[7:4] = 4'd5;
        {2'd2, 4'd14}: S[7:4] = 4'd9;
        {2'd2, 4'd15}: S[7:4] = 4'd2;
        {2'd3, 4'd0}:  S[7:4] = 4'd6;
        {2'd3, 4'd1}:  S[7:4] = 4'd11;
        {2'd3, 4'd2}:  S[7:4] = 4'd13;
        {2'd3, 4'd3}:  S[7:4] = 4'd8;
        {2'd3, 4'd4}:  S[7:4] = 4'd1;
        {2'd3, 4'd5}:  S[7:4] = 4'd4;
        {2'd3, 4'd6}:  S[7:4] = 4'd10;
        {2'd3, 4'd7}:  S[7:4] = 4'd7;
        {2'd3, 4'd8}:  S[7:4] = 4'd9;
        {2'd3, 4'd9}:  S[7:4] = 4'd5;
        {2'd3, 4'd10}: S[7:4] = 4'd0;
        {2'd3, 4'd11}: S[7:4] = 4'd15;
        {2'd3, 4'd12}: S[7:4] = 4'd14;
        {2'd3, 4'd13}: S[7:4] = 4'd2;
        {2'd3, 4'd14}: S[7:4] = 4'd3;
        {2'd3, 4'd15}: S[7:4] = 4'd12;
endcase
end

always_comb
begin
    case ({xor_result[5], xor_result[0], xor_result[4:1]})
        {2'd0, 4'd0}:  S[3:0] = 4'd13;
        {2'd0, 4'd1}:  S[3:0] = 4'd2;
        {2'd0, 4'd2}:  S[3:0] = 4'd8;
        {2'd0, 4'd3}:  S[3:0] = 4'd4;
        {2'd0, 4'd4}:  S[3:0] = 4'd6;
        {2'd0, 4'd5}:  S[3:0] = 4'd15;
        {2'd0, 4'd6}:  S[3:0] = 4'd11;
        {2'd0, 4'd7}:  S[3:0] = 4'd1;
        {2'd0, 4'd8}:  S[3:0] = 4'd10;
        {2'd0, 4'd9}:  S[3:0] = 4'd9;
        {2'd0, 4'd10}: S[3:0] = 4'd3;
        {2'd0, 4'd11}: S[3:0] = 4'd14;
        {2'd0, 4'd12}: S[3:0] = 4'd5;
        {2'd0, 4'd13}: S[3:0] = 4'd0;
        {2'd0, 4'd14}: S[3:0] = 4'd12;
        {2'd0, 4'd15}: S[3:0] = 4'd7;
        {2'd1, 4'd0}:  S[3:0] = 4'd1;
        {2'd1, 4'd1}:  S[3:0] = 4'd15;
        {2'd1, 4'd2}:  S[3:0] = 4'd13;
        {2'd1, 4'd3}:  S[3:0] = 4'd8;
        {2'd1, 4'd4}:  S[3:0] = 4'd10;
        {2'd1, 4'd5}:  S[3:0] = 4'd3;
        {2'd1, 4'd6}:  S[3:0] = 4'd7;
        {2'd1, 4'd7}:  S[3:0] = 4'd4;
        {2'd1, 4'd8}:  S[3:0] = 4'd12;
        {2'd1, 4'd9}:  S[3:0] = 4'd5;
        {2'd1, 4'd10}: S[3:0] = 4'd6;
        {2'd1, 4'd11}: S[3:0] = 4'd11;
        {2'd1, 4'd12}: S[3:0] = 4'd0;
        {2'd1, 4'd13}: S[3:0] = 4'd14;
        {2'd1, 4'd14}: S[3:0] = 4'd9;
        {2'd1, 4'd15}: S[3:0] = 4'd2;
        {2'd2, 4'd0}:  S[3:0] = 4'd7;
        {2'd2, 4'd1}:  S[3:0] = 4'd11;
        {2'd2, 4'd2}:  S[3:0] = 4'd4;
        {2'd2, 4'd3}:  S[3:0] = 4'd1;
        {2'd2, 4'd4}:  S[3:0] = 4'd9;
        {2'd2, 4'd5}:  S[3:0] = 4'd12;
        {2'd2, 4'd6}:  S[3:0] = 4'd14;
        {2'd2, 4'd7}:  S[3:0] = 4'd2;
        {2'd2, 4'd8}:  S[3:0] = 4'd0;
        {2'd2, 4'd9}:  S[3:0] = 4'd6;
        {2'd2, 4'd10}: S[3:0] = 4'd10;
        {2'd2, 4'd11}: S[3:0] = 4'd13;
        {2'd2, 4'd12}: S[3:0] = 4'd15;
        {2'd2, 4'd13}: S[3:0] = 4'd3;
        {2'd2, 4'd14}: S[3:0] = 4'd5;
        {2'd2, 4'd15}: S[3:0] = 4'd8;
        {2'd3, 4'd0}:  S[3:0] = 4'd2;
        {2'd3, 4'd1}:  S[3:0] = 4'd1;
        {2'd3, 4'd2}:  S[3:0] = 4'd14;
        {2'd3, 4'd3}:  S[3:0] = 4'd7;
        {2'd3, 4'd4}:  S[3:0] = 4'd4;
        {2'd3, 4'd5}:  S[3:0] = 4'd10;
        {2'd3, 4'd6}:  S[3:0] = 4'd8;
        {2'd3, 4'd7}:  S[3:0] = 4'd13;
        {2'd3, 4'd8}:  S[3:0] = 4'd15;
        {2'd3, 4'd9}:  S[3:0] = 4'd12;
        {2'd3, 4'd10}: S[3:0] = 4'd9;
        {2'd3, 4'd11}: S[3:0] = 4'd0;
        {2'd3, 4'd12}: S[3:0] = 4'd3;
        {2'd3, 4'd13}: S[3:0] = 4'd5;
        {2'd3, 4'd14}: S[3:0] = 4'd6;
        {2'd3, 4'd15}: S[3:0] = 4'd11;
endcase
end


// P permutation
logic [31:0]P;
assign P = {S[16], S[25], S[12], S[11], S[3],  S[20], S[4],  S[15], 
            S[31], S[17], S[9],  S[6],  S[27], S[14], S[1],  S[22], 
            S[30], S[24], S[8],  S[18], S[0],  S[5],  S[29], S[23], 
            S[13], S[19], S[2],  S[26], S[10], S[21], S[28], S[7]};


// output
assign R_out = P ^ L;

endmodule

